//transaction.sv
class transaction;
  randc bit [3:0] d;
  bit[15:0] o ;

endclass
