interface mux_if();
  logic [7:0] d;
  logic [2:0] sel;
  logic y;
  
endinterface 
  
