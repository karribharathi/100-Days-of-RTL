class transaction;

  rand bit  d;
  rand bit  [2:0]    sel;
  bit    [7:0] y;

  

endclass
