class transaction;
randc bit in1;
randc bit in2;
randc bit cin; 
bit sum;
bit cout;
endclass
