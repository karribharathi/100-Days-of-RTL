//interface
interface dec_if;
  logic [3:0] d;
  logic [15:0] o;

endinterface
