interface demux_if();
  logic  d;
  logic [2:0] sel;
  logic [7:0] y;
  
endinterface 
  
