class transaction;

  rand bit[7:0] d;
  rand bit  [2:0]    sel;
  bit    y;

  

endclass
