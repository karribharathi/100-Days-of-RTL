//interface
interface encoder_if;
  logic [3:0] d;
  logic [1:0] o;

endinterface
