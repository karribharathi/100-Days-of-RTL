//transaction.sv
class transaction;
  randc bit [3:0] d;
  bit [1:0] o ;

endclass
